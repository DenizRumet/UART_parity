module Rx_LAB5_DRF(SCin, SDin, PDout, PDready, ParErr);
input SCin;			// clock input, SDin is valid at the rising clock edge
input SDin;			// serial data input

output [7:0] PDout;	// parallel output
output PDready;		// One-clock-cycle output pulse generated after the last serial data bit is received
output ParErr;

			
assign ParErr = ((SDin == ^SR) && (Counter [3:0] == 4'd8)) ? 1'b0 : 1'b1;

reg [7:0] SR;		// storage unit
reg [3:0] Counter;	// counter
reg SRC;			// storage control


// Data control part
always @(posedge SCin)
begin
	if ( (SDin == 1'b1) && (Counter [3:0] == 4'b0) )	// new serial incoming data 
		SRC <= 1'b1;									// set 1 when data is coming
	else
		if (Counter[3:0] == 4'd7)						// all incoming data is arrived
			SRC <= 1'b0;								// no incoming data
		else
			SRC <= SRC;									// incoming data control is idle
end

// Shift Register Part
always @(posedge SCin)
begin
	if (SRC == 1'b1)									// incoming data state
		begin
			SR [7:1] <= SR[6:0];						//	shift the data stored
			SR [0] <= SDin;								//	store the first data coming
		end
	else
		SR [7:0] <= SR [7:0];							// storage idle
end

// Counter Part to control SDin flow
always @(posedge SCin)
begin
	if (SRC == 1'b0)									// no incoming data
		Counter [3:0] <= 4'b0;							// clear the counter
	else
		Counter [3:0] <= Counter [3:0] + 4'b1;			// increment the counter by 1 when data is coming
end


assign PDout [7:0] = SR [7:0];
assign PDready = (Counter [3:0] == 4'd8) ? 1'b1 : 1'b0;

endmodule
